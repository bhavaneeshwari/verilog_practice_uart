
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 03.01.2026 12:34:27
// Design Name: 
// Module Name: tb_uart
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module tb_uart;
reg clk =0,rst =0;
reg rx =1 ;
reg [7:0] dintx;
reg newd;
wire tx;
wire [7:0] doutrx;
wire donetx;
wire donerx;

uarttop #(1000000,9600) dut (clk,rst,rx,dintx,newd,tx,doutrx,donetx,donerx);
always #5 clk = ~clk;

reg [7:0] rx_data=0,tx_data=0;
initial begin 
rst =1;
repeat(5) @(posedge clk)
rst =0;
for (int i =0;i<10;i++)
begin 
rst =0;
newd=1;
dintx = $random();
wait (tx ==0);
@(posedge dut.tx_ins.uclk);
for (int i =0;i<=7;i++)
begin
@(posedge dut.tx_ins.uclk);
tx_data = {tx,tx_data[7:1]};
end
@(posedge donetx);
end 
for (int i =0;i<=10;i++)
begin 
rst =0;
newd=0;
rx =1'b0;

@(posedge dut.tx_ins.uclk);
for (int i =0;i<=7;i++)
begin
@(posedge dut.tx_ins.uclk);
rx =$random();
rx_data = {rx,rx_data[7:1]};
end
@(posedge donerx);
end 
end 

endmodule
